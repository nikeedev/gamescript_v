module gamescript

struct Vector2
{
mut:
	int x;
	int y;
}

