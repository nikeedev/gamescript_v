module gamescript

pub struct Vector2
{
pub mut:
	x int
	y int
}

